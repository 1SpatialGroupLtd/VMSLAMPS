window pos 100 150
window size 224 125

name console "cmd1_menu"
name parent  "cmd0_menu"

font 0
!8 x 14 pixels
on border
ret code 999

ret text "cmd11_menu"
button text 0 94  " 1 "
ret text "cmd12_menu"
button text 0 80  " 2 "
ret text "cmd13_menu"
button text 0 66  " 3 "
ret text "cmd14_menu"
button text 0 52  " 4 "
ret text "cmd15_menu"
button text 0 38  " 5 "
ret text "cmd16_menu"
button text 0 24  " 6 "

ret text "cmd0_menu"
button text 0  0  "  Exit this Menu            "

