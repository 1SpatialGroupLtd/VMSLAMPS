
!
! E X A M P L E   C D L   F I L E
!
! M E N U  4

! menu placed at lower left of screen
window pos 160 300
window size 120 210

! this is 'menu_4' with a parent menu of 'menu_2'
name console "menu_4"
name parent "menu_2"

!
! Print a title
font 1
add text 0 185 "DIGITISING" 
add text 0 170 "   MENU   "
 
! text is to be output in font 0, and buttons are not to have a border
font 0
off border

! subsequent buttons post text to the mailbox

! this button posts the LITES command 'select all' to the mailbox and
! clears previous selections made by TOGGLE buttons
return code 995
return text "%select all"
button text 0 145  "   SELECT ALL    "

return code 1

! this button posts the LITES command '%select fc 10' to the mailbox
return text "%select fc 10"
toggle text 0 130  "     ROADS       "

! this button posts the LITES command '%select fc 15' to the mailbox
return text "%select fc 15"
toggle text 0 115  "     RIVERS      "

! this button posts the LITES command '%select fc 22' to the mailbox
return text "%select fc 22"
toggle text 0 100  "    CONTOURS     "

! this button posts the LITES command 'start' to the mailbox
offset 0 14
return text "%start"
button text 0 60   "     START       "

! this button posts the LITES command 'end' to the mailbox
return text "%end"
button text 0 45   "      END        "

! this button posts the LITES command 'abandon' to the mailbox
return text "%abandon"
button text 0 30   "    ABANDON      "

! this button causes 'menu_3' to be displayed
on border
return code 993
return text "/%mess exiting/menu_3/"
button text 25 5  " E X I T "
