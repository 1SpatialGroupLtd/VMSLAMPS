window pos 200 100
window size 300 125

name console "cmd15_menu"
name parent  "cmd1_menu"

font 0
!8 x 14 pixels
on border
ret code 1

icon file "up_arrow"
ret text "up"
button icon 10 10
icon file "down_arrow"
ret text "down"
button icon 10 70
icon file "up_arrow"
ret text "up"
button icon 50 10
icon file "down_arrow"
ret text "down"
button icon 50 70
icon file "left_arrow"
ret text "left"
button icon 90 10
icon file "right_arrow"
ret text "right"
button icon 90 70
icon file "inside_box"
ret text "inside"
button icon 130 10
icon file "outside_box"
ret text "outside"
button icon 130 70
icon file "move_box"
ret text "move"
button icon 210 10
icon file "size_box"
ret text "size"
button icon 210 70

