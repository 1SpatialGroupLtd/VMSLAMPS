!! E X A M P L E   C D L   F I L E!! MENU_1 !! menu placed at top centre of screenwindow pos 455 700window size 90 140! this is 'menu_1' with a parent menu of 'cdl$none'name console "menu_1"name parent "cdl$none"! text is to be output in font 0, and buttons are not to have a borderfont 0off border! this button causes UISMENUS to completereturn code 991return text " "button text 0 5  "  S T O P   "return code 999return text "menu_2"button text 0 25  "   LITES2   "! draw a lineadd line 0 45 90 45! define an iconicon file "LSL_LOGO"! this places an icon in the menu (with null ouput)return text "%null"button icon 21 50!add text 0 120 "  Example  "add text 0 105 "   Menus   "