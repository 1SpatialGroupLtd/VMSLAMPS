
!
! E X A M P L E   C D L   F I L E
!
! M E N U  5

! menu placed at lower left of centre of screen
window pos 320 300
window size 120 210

! this is 'menu_5' with a parent menu of 'menu_2'
name console "menu_5"
name parent "menu_2"

!
! Print a title
font 1
add text 0 185 "  EDITING  " 
add text 0 170 "   MENU   "

! subsequent buttons post text to the mailbox
font 0
return code 1

add text 0 140 "     CURSOR     "
! start a group
group
on border

! this button posts the LITES command '%disable big' to the mailbox
return text "%disable big"
choice text 5 125 " SMALL "

! this button posts the LITES command '%enable big' to the mailbox
return text "%enable big"
choice text 75 125 " BIG "

! text is to be output in font 0, and buttons are not to have a border
font 0
off border

! this button posts the LITES command '%zoom 10' to the mailbox
return text "%zoom 10"
button text 0 105  "   ZOOM LOTS      "

! this button posts the LITES command '%zoom 1' to the mailbox
return text "%zoom 1"
button text 0 90   "     CENTRE       "

! this button posts the LITES command '%zoom 0.5' to the mailbox
return text "%zoom 0.5"
button text 0 75   "    ZOOM OUT      "

! this button posts the LITES command '%find' to the mailbox
return text "%find"
button text 0 55   "      FIND         "

! this button posts the LITES command '%delete' to the mailbox
return text "%delete"
button text 0 40   "     DELETE        "

! this button posts the LITES command '%abandon' to the mailbox
return text "%abandon"
button text 0 20   "    ABANDON      "

!
on border
return code 999
return text "menu_3"
button text 25 5  " E X I T "
