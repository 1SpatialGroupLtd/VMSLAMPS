
!
! E X A M P L E   C D L   F I L E
!
! MENU_1 
!

! menu placed at top centre of screen
window pos 455 700
window size 90 140

! this is 'menu_1' with a parent menu of 'cdl$none'
name console "menu_1"
name parent "cdl$none"

! text is to be output in font 0, and buttons are not to have a border
font 0
off border

! this button causes UISMENUS to complete
return code 991
return text " "
button text 0 5  "  S T O P   "

return code 999
return text "menu_2"
button text 0 25  "   LITES2   "

! draw a line
add line 0 45 90 45

! define an icon
icon file "LSL_LOGO"

! this places an icon in the menu (with null ouput)
return text "%null"
button icon 21 50

!
add text 0 120 "  Example  "
add text 0 105 "   Menus   "
