
!
! E X A M P L E   C D L   F I L E
! 
!  M E N U  3
!

! menu placed at middle right of screen
window pos 550 600
window size 90 60
window noframe

! this is 'menu_3' with a parent menu of 'menu_1'
name console "menu_3"
name parent "menu_1"

! text is to be output in font 0, and buttons are not to have a border
font 0
off border

! this button causes the text '%ABAN#%QUIT#%QUIT' to be posted to the mailbox
! and uismenus to complete.
return code 998
return text "%ABAN#%QUIT#%QUIT"
button text 0 10  "  CONFIRM   "

font 1
add text 0 35 " EXIT  "
