window pos 100 150
window size 224 125

name console "cmd0_menu"
name parent  "cdl$none"

font 0
!8 x 14 pixels
off border
ret code 999

ret text "cmd1_menu"
button text 0 84  " 1 "
ret text "cmd2_menu"
button text 0 70  " 2 "
ret text "cmd3_menu"
button text 0 56  " 3 "
ret text "cmd4_menu"
button text 0 42  " 4 "
ret text "cmd5_menu"
button text 0 28  " 5 "
ret text "cmd6_menu"
button text 0 14  " 6 "

