!! E X A M P L E   C D L   F I L E!! M E N U  5! menu placed at lower left of centre of screenwindow pos 320 300window size 120 210! this is 'menu_5' with a parent menu of 'menu_2'name console "menu_5"name parent "menu_2"!! Print a titlefont 1add text 0 185 "  EDITING  " add text 0 170 "   MENU   "! subsequent buttons post text to the mailboxfont 0return code 1add text 0 140 "     CURSOR     "! start a groupgroupon border! this button posts the LITES command '%disable big' to the mailboxreturn text "%disable big"choice text 5 125 " SMALL "! this button posts the LITES command '%enable big' to the mailboxreturn text "%enable big"choice text 75 125 " BIG "! text is to be output in font 0, and buttons are not to have a borderfont 0off border! this button posts the LITES command '%zoom 10' to the mailboxreturn text "%zoom 10"button text 0 105  "   ZOOM LOTS      "! this button posts the LITES command '%zoom 1' to the mailboxreturn text "%zoom 1"button text 0 90   "     CENTRE       "! this button posts the LITES command '%zoom 0.5' to the mailboxreturn text "%zoom 0.5"button text 0 75   "    ZOOM OUT      "! this button posts the LITES command '%find' to the mailboxreturn text "%find"button text 0 55   "      FIND         "! this button posts the LITES command '%delete' to the mailboxreturn text "%delete"button text 0 40   "     DELETE        "! this button posts the LITES command '%abandon' to the mailboxreturn text "%abandon"button text 0 20   "    ABANDON      "!on borderreturn code 999return text "menu_3"button text 25 5  " E X I T "