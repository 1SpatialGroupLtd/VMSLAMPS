window pos 100 150
window size 224 125

name console "cmd2_menu"
name parent  "cmd0_menu"

font 0
!8 x 14 pixels
on border
ret code 999

ret text "cmd21_menu"
button text 0 94  " 1 "
ret text "cmd22_menu"
button text 0 80  " 2 "
ret text "cmd23_menu"
button text 0 66  " 3 "
ret text "cmd24_menu"
button text 0 52  " 4 "
ret text "cmd25_menu"
button text 0 38  " 5 "
ret text "cmd26_menu"
button text 0 24  " 6 "

ret text "cmd0_menu"
button text 0  0  "  Exit this Menu            "

