!! E X A M P L E   C D L   F I L E! !  M E N U  3!! menu placed at middle right of screenwindow pos 550 600window size 90 60window noframe! this is 'menu_3' with a parent menu of 'menu_1'name console "menu_3"name parent "menu_1"! text is to be output in font 0, and buttons are not to have a borderfont 0off border! this button causes the text '%ABAN#%QUIT#%QUIT' to be posted to the mailbox! and uismenus to complete.return code 998return text "%ABAN#%QUIT#%QUIT"button text 0 10  "  CONFIRM   "font 1add text 0 35 " EXIT  "