
!
! E X A M P L E   C D L   F I L E
!
! M E N U 2
!

! menu placed at middle left of screen
window pos 200 495
window size 250 150

! this is 'menu_2' with a parent menu of 'menu_1'
name console "menu_2"
name parent "menu_1"

! text is to be output in font 0, and buttons are to have a border
font 0
on border
!
! this button causes 'menu_4' to be reinitialised and displayed
return code 994
return text "menu_4"
button text 10 30  " DIGITISE "
!
! this button causes 'menu_5' to be reinitialised and displayed
! and the first part of the return text posted to the mailbox
return code 992
return text "/%mess change to editing/menu_5/"
button text 105 30  " EDIT "

! this button causes 'menu_3' to be displayed
return code 999
return text "menu_3"
button text 170 30  " E X I T "
!
! Print a banner
font 2
off border
add text 35 75 " L I T E S"

!
! this button causes 'menu_1' to be displayed
font 0
on border
return code 999
return text "menu_1"
button text 170 130 " RETURN "
