window pos 100 150
window size 224 125

name console "cmd4_menu"
name parent  "cmd0_menu"

font 0
!8 x 14 pixels
on border
ret code 999

ret text "cmd41_menu"
button text 0 94  " 1 "
ret text "cmd42_menu"
button text 0 80  " 2 "
ret text "cmd43_menu"
button text 0 66  " 3 "
ret text "cmd44_menu"
button text 0 52  " 4 "
ret text "cmd45_menu"
button text 0 38  " 5 "
ret text "cmd46_menu"
button text 0 24  " 6 "

ret text "cmd0_menu"
button text 0  0  "  Exit this Menu            "

